../_common/r65c02tc_fsm_intnmi.vhdl