../_common/T65_ALU.vhdl