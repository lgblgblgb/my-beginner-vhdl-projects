../_common/r65c02tc_regbank_axy.vhdl