../_common/T65_Pack.vhdl