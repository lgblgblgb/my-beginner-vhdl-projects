../_common/T65_MCode.vhdl