../_common/T65.vhdl