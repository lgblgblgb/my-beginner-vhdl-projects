../_common/via6522.vhdl