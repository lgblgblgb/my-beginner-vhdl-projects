../_common/r65c02tc_fsm_execution_unit.vhdl