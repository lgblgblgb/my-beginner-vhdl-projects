../_common/r65c02tc_reg_sp.vhdl