../_common/r65c02tc_r65c02_tc_config.vhdl