../_common/r65c02tc_core.vhdl