../_common/r65c02tc_reg_pc.vhdl